/*=========================================================================
===========================================================================
    =            Proyecto:      Práctica 1                            =
    =            Archivo:       compl1.v                              =
    =            Autor:         Adrián Epifanio R.H                   =
    =            Fecha:         08/11/2018                            =
    =            Asignatura:    Estructuras de computadores           =
    =            Lenguaje:      Verilog                               = 
===========================================================================          
=========================================================================*/


/*===================================================================
=                            MODULE                                 =
===================================================================*/
module compl1(output wire [3:0] Sal, input wire [3:0] Ent, input wire cpl);
		
	assign Sal = cpl ? ~Ent : Ent;

endmodule

/*===================================================================*/
/*=========================  End of module  =========================*/
/**
 *
 *
 *   Autor: Adrián Epifanio R.H
 *   Fecha: 08/11/2018
 *
 *
**/

