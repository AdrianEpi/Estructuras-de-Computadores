/*=========================================================================
===========================================================================
    =            Proyecto:      Práctica 1                            =
    =            Archivo:       cl.v                                  =
    =            Autor:         Adrián Epifanio R.H                   =
    =            Fecha:         08/11/2018                            =
    =            Asignatura:    Estructuras de computadores           =
    =            Lenguaje:      Verilog                               = 
===========================================================================          
=========================================================================*/


/*===================================================================
=                            MODULE                                 =
===================================================================*/
module cl(output wire out, input  wire a, b, input wire [1:0] s);

	wire c00, c01, cxor, cnot;
	and	and1(c00, a, b);
	or	or1(c01, a, b);
	xor	puertaxor(cxor, a, b);
	not 	not1(cnot,a);
	
	mux4_1 muliplex1(out, c00, c01, cxor, cnot, s);

endmodule

/*===================================================================*/
/*=========================  End of module  =========================*/
/**
 *
 *
 *   Autor: Adrián Epifanio R.H
 *   Fecha: 08/11/2018
 *
 *
**/

